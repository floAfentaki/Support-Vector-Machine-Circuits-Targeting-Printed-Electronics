parameter N_features = 11,
parameter feature_bits = 4,
parameter weightWidth = 6,
parameter  biasWidth= 6,
parameter  inputWidth= 4,
parameter [weightWidth*N_features-1: 0] weights[0 : 20]= {66'b000001000000000000000001000100000010000011000011111110111111110110, 66'b000111001001000011111010000100000110000010111111000010111110111000, 66'b000111001000111111111100000110001001111111111111000001111110111011, 66'b000011000010111111111111000001000101111111111111000001111111111111, 66'b000100000000111111000000000001000110111111111110000001000000000001, 66'b000101111011111111000100000101001010000001000000000001111101000011, 66'b111101000011111110111110000100111100000000000010111100000010111000, 66'b000100010110000101101000000010101010111111000000111101000001101010, 66'b000111011101000011100111001000101100111010000011111101111110101101, 66'b000110010000111110110010111110110001111101000101000001111111111001, 66'b000101001010000000111001111111111000111100000100000011000000000001, 66'b111101000001111111111111000100111111000001000010111101000001111100, 66'b000011001011000010110000000000110001000011001000000000111110101010, 66'b000001011000000000101100001010111010000000010001111101111011101000, 66'b000011010001000000110011000000111000000011000111111110111101110000, 66'b111110000000000000000000000100111111000001000010111110000000111111, 66'b111111000010000011111000000001110110000010000110111110000000111001, 66'b111101000110000011110011001100111100000000010001111100111101110111, 66'b111101000000111111000000000011000000000001000001111110000001000000, 66'b000000000001000010111001111000110100000010000000000000000001111100, 66'b111011000000111110000001000100000000000011000001111101000001111111 },
parameter [weightWidth-1 : 0] bias[0 : 20]= {6'b000111, 6'b111001, 6'b110111, 6'b110111, 6'b110110, 6'b110111, 6'b001100, 6'b000111, 6'b000001, 6'b111011, 6'b110111, 6'b001011, 6'b001101, 6'b001000, 6'b000010, 6'b001001, 6'b001011, 6'b001000, 6'b001001, 6'b001000, 6'b001001 }