parameter N_features = 33,
parameter feature_bits = 6,
parameter weightWidth = 4,
parameter  biasWidth= 4,
parameter  inputWidth= 4,
parameter [weightWidth*N_features-1: 0] weights[0 : 14]= {132'b000000010001000000010000101100001111000011110000000000100000000000000000000100110011010000010010000000010000111000001110110000010000, 132'b000100010011110100100000000000000010000100010000000001001001000011100000000101000000010100100010000000010000111100000000000011110000, 132'b000100010001001011110000000000000010001000010000000000110000110100000000000001000110010100100000000000000000110011110000000000000000, 132'b000000010000000000001110000011100001000100001111000000100000111100000000000000100010001000010000111000001111111111100000000000001110, 132'b000000000010111100110000000000000011000100000000111000000000110100000000000001010100010100000001000000000000100100000000000000000000, 132'b000000000001000100000000100100001101111111100000000100110000001000000000000011110000000000000000000000000000001100001100100100000000, 132'b000000100010000000000000111100000000000000000000010001001001001111101101000000001010000000000000000000000000011000000000000000001111, 132'b001001100000011010010000000100000100000100010000011001100000110100101110110100000000000000110000000010010000010000000000000011000010, 132'b000000100000000011111100000011100000000000001110000000011111000100001111000000000000000000001111110111111110000111010000000000001110, 132'b000011110000000100000010110100011110111111110001000000000000000100000000000000000000000000000000001000000001000000101111111000000010, 132'b111111110000000000010100111100100000000000000001000000001101000111111111000000001110000000000001001000010010000100110000000000000011, 132'b000011110000001011100100000000110000000000000010000011110001000000000000000000000000000000000001001100000010000000110000000000000100, 132'b000000000001000000100000100100001101111111100000000000010000001000001111000100000000000000000000000000010000000000001100101000100000, 132'b000000000100110001000000111100000000000000000000000000011001001111110000001000001010000000000000000000100000010000000000000000011111, 132'b000000001111001000000000110100001101111011010000000000000101000100010001111111110011000000000000000000000000111000001101101100010000 },
parameter [weightWidth-1 : 0] bias[0 : 14]= {4'b1111, 4'b1110, 4'b1011, 4'b0000, 4'b1110, 4'b0001, 4'b0000, 4'b1100, 4'b0100, 4'b1111, 4'b1110, 4'b1100, 4'b0011, 4'b0001, 4'b0001 }