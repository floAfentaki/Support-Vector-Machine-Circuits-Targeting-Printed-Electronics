parameter N_features = 11,
parameter feature_bits = 4,
parameter weightWidth = 5,
parameter  biasWidth= 5,
parameter  inputWidth= 4,
parameter [weightWidth*N_features-1: 0] weights[0 : 20]= {55'b0000000000000000000100011000010001100010111111111110110, 55'b0011101001000101101000100001100000100000000011111011000, 55'b0011000111000001110000110010011111111111000001111011100, 55'b0001100001000001111100001001000000011111000000000000000, 55'b0010000000000000000000001001011111111111000010000000000, 55'b0010111100000000010000101010100000100000000011111000010, 55'b1111000011111111111100100111010000000001111000001011000, 55'b0001101110001011000100001100011111100000111010000110001, 55'b0011101110000111000101000100011101100010111101111010001, 55'b0011001110111111001111111100101110100101000001111111001, 55'b0010001010000001100111111110011110000100000100000000001, 55'b1111000000111111111100100111110000000010111100000011101, 55'b0001001011000011000100000100100001100111000001111010001, 55'b0000101110000001000101001110100000001110111101101110001, 55'b0001001110000001001100000110010001100110111111110110001, 55'b1111000000000000000000011000000000000001111110000000000, 55'b0000000001000101100100001101110000100101111110000011010, 55'b1111000110000101010001100111000000001110111001111010111, 55'b1111000000111110000000011000000000100001111110000000000, 55'b0000000000000101100111001101000001000000000000000111100, 55'b1101100000111110000000011000000001000001111100000100000 },
parameter [weightWidth-1 : 0] bias[0 : 20]= {5'b00111, 5'b11001, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b01100, 5'b00111, 5'b00000, 5'b11011, 5'b10111, 5'b01011, 5'b01100, 5'b01000, 5'b00010, 5'b01001, 5'b01010, 5'b00111, 5'b01001, 5'b01000, 5'b01001 }
