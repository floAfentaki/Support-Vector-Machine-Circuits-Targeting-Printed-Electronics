parameter N_features = 33,
parameter feature_bits = 6,
parameter weightWidth = 5,
parameter  biasWidth= 5,
parameter  inputWidth= 4,
parameter [weightWidth*N_features-1: 0] weights[0 : 14]= {165'b000000001000011000000001000000101010000011101000001111000000000000010000000000001111111111000110011000110010010001000100000000001100000111000000011011110000001000000, 165'b000100001100111110100010100000111110000000100000110001100000000000100010010111111110000000000100100000000010110010000100000000001100000111010000011111000001111000000, 165'b000100001000010001001110100000000000000000101001010001000000000000011000000110101111100000000000100101100010100010100001000000000100000101111110100000000000000000000, 165'b000010001100000000000000111011000001110000011000100000111101000000010011111111100000000000000010010000101001000001000000111000000011101111011110000000000000000011011, 165'b000000000100101111100011000000000000000000111000110000100000111001111100000110011111100001000010101001000010110000000011000000000100000100010000000000000000000100000, 165'b000010000000010000100000000000100010000011001111011101100000000110011000000001010000011111000001111011111000000000000000000000000000000001100000010111100100000100001, 165'b000000010000100000000000000000111100000000000000000000000000010000100010001001111101111001000010000010100111110000100000000000000000000011010000011111000000000011110, 165'b001000110000001011001000100000000110000001000000100001000000011010111000000110100010111100110100000000000000000011100000000001000100000010010000000000000001011100101, 165'b000000010111111111111111010111000001101100000000000000011011000010001111110000110000011110111110000000000000000000011101110011111011011000111100100000000000000011011, 165'b111111111000001000100000100101110100001111100111101111000011000011111100001000100000011111000000000000000000000000000001001000000100011000000010011110110110000000100, 165'b111101111000001111110001001000111100010100000000000000000011000000000011010000101111011110000010000011100000000000000011001000001000100000110011000000000000000000110, 165'b111111111000000001001110001001000000011000000000010000000100000011111000011111110000000000111110000000000000000000000011001100000000100111110011000000000000000001001, 165'b000001111100011111110010000000100100000011001111011101100000000000001000000001000000011110000101111111111000000000000000000000001100000000010000011000100110010011111, 165'b000001111101000110000100100000111010000000000000000000000000000010001010001001101111011111001010000010011111110000000000000000010000000010000000011111000000001011110, 165'b111110000011110001010000000000110100000011001110111101000000000001111101011000100001100011111101111000110000010000000000000000000000000110110000011010101010001000000 },
parameter [weightWidth-1 : 0] bias[0 : 14]= {5'b11110, 5'b11100, 5'b10110, 5'b00001, 5'b11011, 5'b00011, 5'b00000, 5'b11000, 5'b01000, 5'b11101, 5'b11011, 5'b10111, 5'b00110, 5'b00010, 5'b00010 }
