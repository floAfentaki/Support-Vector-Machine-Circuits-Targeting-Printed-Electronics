parameter N_features = 11,
parameter feature_bits = 4,
parameter weightWidth = 6,
parameter  biasWidth= 6,
parameter  inputWidth= 4,
parameter [weightWidth*N_features-1: 0] weights[0 : 14]= {66'b111111010001110100000000001001000011111110010000001001111000100011, 66'b111111011110000000111101001100000000111100000110000101110011100101, 66'b000101010111000010000000001100000000110010000010001000110100110100, 66'b000100001111000011000010000111000001110011000000000111111100111011, 66'b000111010001000010000011001010111101111001001001000011111010110111, 66'b111000001100110100001101010010111110000010001111010001110011100001, 66'b110111011110000010001010010101111001000101111010001010100110100001, 66'b000110010101000100001011001101111010110101110010001100110100110001, 66'b000110001011000011001110000101111110110011110010001011000000111101, 66'b000111000110110000000100001010000001001011010001001110110010100010, 66'b110010011101111100110010010010111010011010010011111101100001100001, 66'b111011010101000011111000001111110110011110000101111110100110100100, 66'b000001111101111100111011001010000001000101000110001001110100101111, 66'b110001010010111111101110001101000110001000001111111110100111101100, 66'b000001110111111110000010000111111110000100000101001011111100110011 },
parameter [weightWidth-1 : 0] bias[0 : 14]= {6'b111101, 6'b110001, 6'b101000, 6'b101000, 6'b101010, 6'b001000, 6'b000001, 6'b110001, 6'b101111, 6'b001101, 6'b001101, 6'b000011, 6'b010011, 6'b001111, 6'b001111 }